module GenRoundKeys(K0, K1, K2, K3, K4, K5, K6, K7, K8, K9, K10);
	input [127:0] K0;
	output [127:0] K1, K2, K3, K4, K5, K6, K7, K8, K9, K10;
	wire [31:0] rcon0, rcon1, rcon2, rcon3, rcon4, rcon5, rcon6, rcon7, rcon8, rcon9, rcon10;
	wire [31:0] w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43;
	wire [31:0] rw3, rw7, rw11, rw15, rw19, rw23, rw27, rw31, rw35, rw39;
	wire [31:0] sw3, sw7, sw11, sw15, sw19, sw23, sw27, sw31, sw35, sw39;
	
	assign rcon1  = 32'h01000000;
	assign rcon2  = 32'h02000000;
	assign rcon3  = 32'h04000000;
	assign rcon4  = 32'h08000000;
	assign rcon5  = 32'h10000000;
	assign rcon6  = 32'h20000000;
	assign rcon7  = 32'h40000000;
	assign rcon8  = 32'h80000000;
	assign rcon9  = 32'h1b000000;
	assign rcon10 = 32'h36000000;

	assign {w0,w1,w2,w3} = K0;
	assign K1 = {w4,w5,w6,w7};
	assign K2 = {w8,w9,w10,w11};
	assign K3 = {w12,w13,w14,w15};
	assign K4 = {w16,w17,w18,w19};
	assign K5 = {w20,w21,w22,w23};
	assign K6 = {w24,w25,w26,w27};
	assign K7 = {w28,w29,w30,w31};
	assign K8 = {w32,w33,w34,w35};
	assign K9 = {w36,w37,w38,w39};
	assign K10 = {w40,w41,w42,w43};

	RotWord R0(w3, rw3);
	SubWord S0(rw3, sw3);
	assign w4 = w0^sw3^rcon1;
	assign w5 = w4^w1;
	assign w6 = w5^w2;
	assign w7 = w6^w3;
	RotWord R1(w7, rw7);
	SubWord S1(rw7, sw7);
	assign w8 = w4^sw7^rcon2;
	assign w9 = w8^w5;
	assign w10 = w9^w6;
	assign w11 = w10^w7;
	RotWord R2(w11, rw11);
	SubWord S2(rw11, sw11);
	assign w12 = w8^sw11^rcon3;
	assign w13 = w12^w9;
	assign w14 = w13^w10;
	assign w15 = w14^w11;
	RotWord R3(w15, rw15);
	SubWord S3(rw15, sw15);
	assign w16 = w12^sw15^rcon4;
	assign w17 = w16^w13;
	assign w18 = w17^w14;
	assign w19 = w18^w15;
	RotWord R4(w19, rw19);
	SubWord S4(rw19, sw19);
	assign w20 = w16^sw19^rcon5;
	assign w21 = w20^w17;
	assign w22 = w21^w18;
	assign w23 = w22^w19;
	RotWord R5(w23, rw23);
	SubWord S5(rw23, sw23);
	assign w24 = w20^sw23^rcon6;
	assign w25 = w24^w21;
	assign w26 = w25^w22;
	assign w27 = w26^w23;
	RotWord R6(w27, rw27);
	SubWord S6(rw27, sw27);
	assign w28 = w24^sw27^rcon7;
	assign w29 = w28^w25;
	assign w30 = w29^w26;
	assign w31 = w30^w27;
	RotWord R7(w31, rw31);
	SubWord S7(rw31, sw31);
	assign w32 = w28^sw31^rcon8;
	assign w33 = w32^w29;
	assign w34 = w33^w30;
	assign w35 = w34^w31;
	RotWord R8(w35, rw35);
	SubWord S8(rw35, sw35);
	assign w36 = w32^sw35^rcon9;
	assign w37 = w36^w33;
	assign w38 = w37^w34;
	assign w39 = w38^w35;
	RotWord R9(w39, rw39);
	SubWord S9(rw39, sw39);
	assign w40 = w36^sw39^rcon10;
	assign w41 = w40^w37;
	assign w42 = w41^w38;
	assign w43 = w42^w39;
endmodule
