`timescale 1 ns / 100 ps
module MixColumns_tb;
	integer a;
	reg [127:0] i = 128'hdb13534500000000f20a225c;
	wire [127:0] o;
	MixColumns M(i, o);
	initial begin
		#1;
		$display("i:%h, o:%h", i, o);
		$finish;
	end
endmodule
